module SpectralShaper (
    input clk_x25,
    input [7:0] i_I,
    input [7:0] i_Q,
    
);




endmodule
